# Svenska str�ngar skrivna av Sebastian Rasmussen.

0.0:  FDTUI �r ett TUI-skal f�r FreeDOS.
0.1:  Copyright (C) 2017-2021 Ercan Ersoy
0.2:  FDTUI licensierat under GNU GPL version 2 och GNU GPL version 3.

1.0:Kan inte initiera FDOSTUI-subsystemet.
1.1:\r\nTryck p� valfri tangent f�r att �terg� till DOSSHELL.

2.0:Interna program
2.1:Filhanterare
2.2:K�r

3.0:Avsluta
3.1:Avsluta

4.0:Filhanterare

5.0:Arkiv
5.1:�ppna
5.2:Ny katalog
5.3:Avsluta

6.0:Redigera
6.1:Klipp ut
6.2:Kopiera
6.3:Klistra in
6.4:Byt namn
6.5:�ndra attribut
6.6:Arkiv
6.7:G�md
6.8:Skrivskyddad
6.9:System
6.10:Ta bort

7.0:Visa
7.1:Uppdatera
7.2:Visa arkivobjekt
7.3:Visa g�mda objekt
7.4:Visa skrivskyddade objekt
7.5:Visa systemobjekt

8.0:G�
8.1:Bak�t
8.2:Fram�t
8.3:Upp

9.0:Ny katalog
9.1:Katalognamn:

10.0:Byt namn
10.1:Nytt namn:

11.0:Objektattribut:

12.0:K�r
12.1:Kommando att k�ra:
